`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Southern Methodist University
// Engineer: Wei Zhang
// 
// Create Date: 09/30/2020 02:37:48 PM
// Design Name: simple_readout_bt.v
// Module Name: simple_readout_tb
// Project Name: ETROC1 Array
// Target Devices: KC705
// Tool Versions: Vivado 2018.2
// Description: test bench to simulate simple readout module
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module simple_readout_tb();
reg clock;
reg reset;
reg start;
reg [15:0] write_num;
wire BC0_OUTP;
wire BC0_OUTN;
wire L1ACC_OUTP;
wire L1ACC_OUTN;


initial begin
reset = 1'b0;
clock = 1'b0;
start = 1'b0;
write_num = 16'd12;
#1000 reset = 1'b1;
#100  reset = 1'b0;
#100  start = 1'b0;
#500  start = 1'b1;
#60   start = 1'b0;

#5000000 $stop;
end

always begin
#5 clock = ~clock;
end

simple_readout simple_readout_inst(
.clock(clock),                   // input clock 100 MHz
.reset(reset),                   // reset signal, low active
.start(start),                   // start signal is used to trigger BC0 and L1ACC, generated by config_reg
.write_num(write_num),           // write BC0 and L1ACC loop number
.BC0_OUTP(BC0_OUTP),             // Binary counter clear signal Positive
.BC0_OUTN(BC0_OUTN),             // Binary counter clear signal Negative
.L1ACC_OUTP(L1ACC_OUTP),         // L1 accumulation signal Positive
.L1ACC_OUTN(L1ACC_OUTN)          // L1 accumulation signal Negative
);
endmodule
