`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Southern Modist University
// Engineer: Wei Zhang
// 
// Create Date: 09/30/2020 10:07:08 AM
// Design Name: kc705_mig
// Module Name: simple_readout
// Project Name: ETROC1 Array
// Target Devices: KC705 EVB Board
// Tool Versions: Vivado 2018.2
// Description: 
// 
// Dependencies: 
// 
// Revision: V1.0
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module simple_readout(
input clock,                    // input clock 100 MHz
input reset,                    // reset signal, low active
input start,                    // start signal is used to trigger BC0 and L1ACC, generated by config_reg
input [15:0] write_num,          // write BC0 and L1ACC loop number
output BC0_OUTP,                // Binary counter clear signal Positive
output BC0_OUTN,                // Binary counter clear signal Negative
output L1ACC_OUTP,              // L1 accumulation signal Positive
output L1ACC_OUTN               // L1 accumulation signal Negative
);
reg BC0;
reg L1ACC;
reg [15:0] write_reg;
reg [10:0] counter_reg;
always @(posedge clock)
begin
    if(reset)
        counter_reg <= 1'b0;
    else
        if(start)
            counter_reg <= 1'b0;
        else
            counter_reg <= counter_reg + 1'b1;
end;

reg [13:0] delay_num;
// state machine define
reg [2:0] current_state, next_state;
localparam state_inital = 3'd0;
localparam state_1 = 3'd1;
localparam state_2 = 3'd2;
localparam state_3 = 3'd3;
localparam state_4 = 3'd4;
localparam state_5 = 3'd5;
localparam state_6 = 3'd6;

always @(posedge clock)
begin
    if(reset)
        current_state <= state_inital;      // reset to state_inital  
    else
        current_state <= next_state;        // move to next state
end

reg [10:0]Counter_V;

always @(posedge clock)
begin
    if(reset)                                   // reset to initial state 
    begin
        next_state <= state_inital;
        delay_num <= 13'd0;
    end
    else
    begin
        case(current_state)
        state_inital:                           // initial state
            begin
                BC0 <= 1'b0;                    // initial BC0 to low
                L1ACC <= 1'b0;                  // initial L1ACC to low
                if(start)                       // start signal enable or disable state machine
                begin
                    write_reg <= write_num;
                    next_state <= state_1;
                end
                else
                    next_state <= state_inital;
            end
        state_1:                                            // state_1
            if(write_reg != 0)
            begin
                Counter_V <= counter_reg;
                write_reg <= write_reg - 1'b1; 
                next_state <= state_2;    
            end
            else
                next_state <= state_inital;
        state_2:
            begin
                if(counter_reg == Counter_V + 10'd100)         //delay 1000 * clock period to assert BC0 to high
                begin
                    BC0 <= 1'b1;
                    Counter_V <= counter_reg;                   // record current counter value
                    next_state <= state_3;                      // move to state_3
                end
                else
                    next_state <= state_2;                      // loop back to state_2
            end 
        state_3:
            begin
                if(counter_reg == Counter_V + 4'd6)             // BC0 signal keep 5*10 ns high
                begin
                    BC0 <= 1'b0;                                // set BC0 = 0
                    Counter_V <= counter_reg;                   // record current counter value
                    next_state <= state_4;                      // move to state_4
                end 
                else
                    next_state <= state_3;                      // loop back to state_3
            end      
        state_4:
            begin
                if(counter_reg == Counter_V + 10'd100)
                begin
                    L1ACC <= 1'b1;                              // set L1ACC = 1
                    Counter_V <= counter_reg;                   // record current counter value
                    next_state <= state_5;                      // move to state_5
                end
                else
                    next_state <= state_4;                      // loop back to state_4
            end
        state_5:
            begin
                if(counter_reg == Counter_V + 4'd6)            
                begin   
                    L1ACC <= 1'b0;                              // set L1ACC = 0
                    delay_num <= 1'b0;
                    next_state <= state_6;                      // loop back to state_6
                end      
                else
                    next_state <= state_5;                      // loop back to state_5
            end 
        state_6:
            begin
                delay_num <= delay_num + 1'b1;
                if(delay_num == 13'd5500)                       // between each frame should have enough time interval
                begin
                    if(write_reg == 0)
                        next_state <= state_inital;             // back to state_inital
                    else
                        next_state <= state_1;                  // back to state_1
                end
                else
                    next_state <= state_6;                      // loop back to state_5
            end   
        endcase
        
    end
end
/*******************************************************************/
// BC0 single-ended to differential
OBUFDS #(
      .IOSTANDARD("LVDS18"),    // Specify the output I/O standard
      .SLEW("SLOW")             // Specify the output slew rate
   ) OBUFDS_BC0_inst(
      .O(BC0_OUTP),             // Diff_p output (connect directly to top-level port)
      .OB(BC0_OUTN),            // Diff_n output (connect directly to top-level port)
      .I(BC0)                   // Buffer input 
   );
/*******************************************************************/
// L1ACC single-ended to differential
OBUFDS #(
      .IOSTANDARD("LVDS18"),    // Specify the output I/O standard
      .SLEW("SLOW")             // Specify the output slew rate
   ) OBUFDS_L1ACC_inst(
      .O(L1ACC_OUTP),           // Diff_p output (connect directly to top-level port)
      .OB(L1ACC_OUTN),          // Diff_n output (connect directly to top-level port)
      .I(L1ACC)                 // Buffer input 
   );
endmodule
